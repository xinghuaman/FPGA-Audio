localparam signed a0 =     0;
localparam signed a1 =   -70;
localparam signed a2 =  -145;
localparam signed a3 =  -226;
localparam signed a4 =  -317;
localparam signed a5 =  -419;
localparam signed a6 =  -535;
localparam signed a7 =  -666;
localparam signed a8 =  -813;
localparam signed a9 =  -977;
localparam signed a10 = -1157;
localparam signed a11 = -1354;
localparam signed a12 = -1566;
localparam signed a13 = -1791;
localparam signed a14 = -2024;
localparam signed a15 = -2264;
localparam signed a16 = -2503;
localparam signed a17 = -2738;
localparam signed a18 = -2961;
localparam signed a19 = -3165;
localparam signed a20 = -3342;
localparam signed a21 = -3484;
localparam signed a22 = -3580;
localparam signed a23 = -3622;
localparam signed a24 = -3601;
localparam signed a25 = -3505;
localparam signed a26 = -3326;
localparam signed a27 = -3053;
localparam signed a28 = -2678;
localparam signed a29 = -2193;
localparam signed a30 = -1589;
localparam signed a31 =  -860;
localparam signed a32 =     0;
localparam signed a33 =   995;
localparam signed a34 =  2129;
localparam signed a35 =  3403;
localparam signed a36 =  4816;
localparam signed a37 =  6368;
localparam signed a38 =  8054;
localparam signed a39 =  9869;
localparam signed a40 = 11806;
localparam signed a41 = 13855;
localparam signed a42 = 16007;
localparam signed a43 = 18249;
localparam signed a44 = 20566;
localparam signed a45 = 22943;
localparam signed a46 = 25364;
localparam signed a47 = 27810;
localparam signed a48 = 30263;
localparam signed a49 = 32703;
localparam signed a50 = 35111;
localparam signed a51 = 37464;
localparam signed a52 = 39744;
localparam signed a53 = 41930;
localparam signed a54 = 44002;
localparam signed a55 = 45942;
localparam signed a56 = 47731;
localparam signed a57 = 49352;
localparam signed a58 = 50791;
localparam signed a59 = 52032;
localparam signed a60 = 53065;
localparam signed a61 = 53879;
localparam signed a62 = 54466;
localparam signed a63 = 54821;
localparam signed a64 = 54939;
